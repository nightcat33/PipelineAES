library verilog;
use verilog.vl_types.all;
entity test_bench_top is
end test_bench_top;
